architecture rtl of I2S_deserializer is
begin
end rtl;
